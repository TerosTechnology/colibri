  constant a : integer := ;
  constant b : unsigned := ;
  constant c : signed := ;
  constant d : std_logic := ;
  constant e : std_logic_vector := ;
  constant f : std_logic_vector(5 downto 0) := ;
  signal g : std_logic;
  signal h : std_logic;
  signal i : std_logic;
