module nonansimodule (  );
  parameter ADDR_WIDTH = 8;              //! Address-bus width.

  reg stop_flag;

endmodule
